library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

ENTITY processor IS
    PORT (
        clock       : in std_logic;
        reset       : in std_logic;
    );
END ENTITY;

ARCHITECTURE processor_arch OF processor IS

BEGIN

END processor_arch;
